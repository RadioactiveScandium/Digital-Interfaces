package top_pkg;

`define DSIZE 4

endpackage